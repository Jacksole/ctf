BZh91AY&SY �f�  �_�Px����߰����PX�&d{Y�HS4���i�����$�@!�h=5SM5 i� ��@�@4��L��byG�#j4 A������&L�20�&�db``D���j<��P��h4  aD�	���J>��-����BEX�#UiU�5����/����_���-qO��<�5$����yfb2*5�p�E��4$�11���x��N�l�Ǧ��O�gK�;B3n�����߃�Щ���ۑ)hn,,e�C�N�eF�fR�S����o��e���z���6�����q#Z�����Z�I���x)%."�t��i��A��T�c8� ��]�B!OKy��%��Y���O��Ը���`���D(���C�M��*��rlV�D����/p�^޵�^�����5���//��ߦ�O��b�)��mv�y���i���M�=7��[
+�<��4u�n<�s�H{��^�=�鬨�M��	�\b�&u�T7]\�#��N#J��sg�6���X���)�q����E5�a�е9IEH*���ܠ5o�L�r*��K.�ūyA}��Em�s]����x�o�}^1������.t�fǺ�	�[���\m��!M��iE��i���<�Po���z%Q�鹲�x�N`�y�Z�9�� �yl`1LYZ-�z��X��ɞr8S�Pz��US)�Qc�ͻ��a�T�X��:5l�9P��f���ey6��-;�T P3܀����Ӡ����f��W�Hl��cͩ���[0��ge�!B}@�x�R�:��m�@���ڂ�S��i�uלb̎���Σ3^f�%q���"�(H R3H�